`ifndef ${t_uvc_name_upper}_SEQ_LIST_SV
`define ${t_uvc_name_upper}_SEQ_LIST_SV

`include "${t_uvc_name}_seq_base.sv"
`include "${t_uvc_name}_random_seq.sv"
`include "${t_uvc_name}_direct_seq.sv"

`endif // ${t_uvc_name_upper}_SEQ_LIST_SV

